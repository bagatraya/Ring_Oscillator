magic
tech sky130A
magscale 1 2
timestamp 1729053058
<< metal1 >>
rect 714 2126 748 2158
rect 165 1847 175 1899
rect 227 1847 237 1899
rect 267 1854 543 1891
rect 583 1854 859 1891
rect 889 1847 899 1899
rect 951 1847 961 1899
rect 100 1616 130 1654
<< via1 >>
rect 175 1847 227 1899
rect 899 1847 951 1899
<< metal2 >>
rect 175 1899 227 1909
rect 899 1899 951 1909
rect 227 1847 899 1899
rect 175 1837 227 1847
rect 899 1837 951 1847
use inverter_gate  x1
timestamp 1729045033
transform 1 0 53 0 1 1306
box -55 9 368 1136
use inverter_gate  x2
timestamp 1729045033
transform 1 0 369 0 1 1306
box -55 9 368 1136
use inverter_gate  x3
timestamp 1729045033
transform 1 0 685 0 1 1306
box -55 9 368 1136
<< labels >>
flabel metal2 874 1870 874 1870 0 FreeSans 160 0 0 0 out
port 0 nsew
flabel metal1 732 2140 732 2140 0 FreeSans 160 0 0 0 vdd
port 1 nsew
flabel metal1 120 1636 120 1636 0 FreeSans 160 0 0 0 gnd
port 2 nsew
<< end >>
